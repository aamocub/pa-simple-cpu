module control_unit #(
    parameter integer DATAWIDTH = 32
) ();

    // TODO: Lista de problemas a tener en cuenta
    // 1. Control de muxes en funcion de opcode

endmodule
