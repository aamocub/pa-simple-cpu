
// Instruction Encoding - 32-bits
// ________________________________________________________________
// | offset[31:19] | ra[18:14] | rb[13:9] | rd[8:4] | opcode[3:0] |
// ----------------------------------------------------------------

module decoder
    import pa_pkg::*;
    import riscv_pkg::*;
(
    input  logic [ 31:0] instr_i,
    output wire  [31:19] offset_o,
    output wire  [18:14] ra_o,
    output wire  [ 13:9] rb_o,
    output wire  [  8:4] rd_o,
    output wire  [  3:0] opcode_o,
    output wire          exception_o
);

endmodule
