// This package includes all parameters, types, enums and others that are required by risc-v.

package riscv_pkg;

    localparam XLEN = 32;

endpackage
