// This package includes all parameters, types, enums and others that are required by the processor itself.

package pa;
endpackage
