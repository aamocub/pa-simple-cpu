/*
    NOTE: The overview of the CPU core. Each stage is divided in its own module. Each module will have a series of inputs and outputs. For the pipeline registers, it will be its own registers, outside of the module. The semi-finished IF stage is an example of this.
*/

module top
    import pa_pkg::*;
    import riscv_pkg::*;
#(
    parameter DEBUG = 0
) (
    input logic clk_i,
    input logic rst_i
);


    // ----------------------------------------------------------------------------------------------------------------
    // IF Stage
    // ----------------------------------------------------------------------------------------------------------------

    // ----------------------------------------------------------------------------------------------------------------
    // ID Stage
    // ----------------------------------------------------------------------------------------------------------------

    // ----------------------------------------------------------------------------------------------------------------
    // EX Stage
    // ----------------------------------------------------------------------------------------------------------------

    // ----------------------------------------------------------------------------------------------------------------
    // M Stage
    // ----------------------------------------------------------------------------------------------------------------

    // ----------------------------------------------------------------------------------------------------------------
    // WB Stage
    // ----------------------------------------------------------------------------------------------------------------


endmodule
