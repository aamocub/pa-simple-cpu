module control_unit #(
    parameter integer DATAWIDTH = 32
) ();

endmodule
