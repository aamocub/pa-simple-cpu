// This package includes all parameters, types, enums and others that are required by risc-v.

package riscv;
endpackage
